class sr_coverage extends uvm_subscriber #(sr_sequence_item);

  //----------------------------------------------------------------------------
  `uvm_component_utils(sr_coverage)

  sr_sequence_item txn;
  real cov;
 
  covergroup dut_cov;
    option.per_instance= 1;
    option.comment     = "dut_cov";
    option.name        = "dut_cov";
    option.auto_bin_max= 4;
    
    S:coverpoint txn.s { 
        bins s_high={1};
        bins s_low ={0};
    }

    R:coverpoint txn.r { 
        bins r_high={1};
        bins r_low ={0};
    }

    SXR:cross S,R;
  endgroup:dut_cov;

function new(string name="sr_coverage",uvm_component parent);
    super.new(name,parent);
    dut_cov=new();
  endfunction

  //---------------------  write method ----------------------------------------
  function void write(sr_sequence_item t);
    txn=t;
    dut_cov.sample();
  endfunction
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  function void extract_phase(uvm_phase phase);
    super.extract_phase(phase);
    cov=dut_cov.get_coverage();
  endfunction
  //----------------------------------------------------------------------------


  //----------------------------------------------------------------------------
  function void report_phase(uvm_phase phase);
    super.report_phase(phase);
    `uvm_info(get_type_name(),$sformatf("Coverage is %f",cov),UVM_MEDIUM)
  endfunction
  //----------------------------------------------------------------------------
  
endclass:sr_coverage
